module hello;
  initial 
    begin
      $display("Hello, bonjour, yo, hi, hola!");
      $finish;
    end
endmodule
